LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY NOTASMUSICALES IS
PORT( CLK, LA, DO, MI, SOL, RE, FA, SI : IN STD_LOGIC;
      SONIDO : OUT STD_LOGIC);
END NOTASMUSICALES;

ARCHITECTURE BEHAVIORAL OF NOTASMUSICALES IS 
--------------------- FRECUENCIAS DE LAS NOTAS ------------------------------
SIGNAL CONT : STD_LOGIC_VECTOR (16 DOWNTO 0) := (OTHERS => '0');
CONSTANT CONT_MAX: STD_LOGIC_VECTOR := "11011101111100100"; --113636(DEC)

SIGNAL CONT1 : STD_LOGIC_VECTOR (17 DOWNTO 0) := (OTHERS => '0');
CONSTANT CONT_MAX1: STD_LOGIC_VECTOR := "101110110001010010"; --191570(DEC)

SIGNAL CONT2 : STD_LOGIC_VECTOR (17 DOWNTO 0) := (OTHERS => '0');
CONSTANT CONT_MAX2: STD_LOGIC_VECTOR := "100101000110100111"; --151975(DEC)

SIGNAL CONT3 : STD_LOGIC_VECTOR (16 DOWNTO 0) := (OTHERS => '0');
CONSTANT CONT_MAX3: STD_LOGIC_VECTOR := "11111001000111111"; --127551(DEC)

SIGNAL CONT4 : STD_LOGIC_VECTOR (17 DOWNTO 0) := (OTHERS => '0');
CONSTANT CONT_MAX4: STD_LOGIC_VECTOR := "101001100100011001"; --170265(DEC)

SIGNAL CONT5 : STD_LOGIC_VECTOR (17 DOWNTO 0) := (OTHERS => '0');
CONSTANT CONT_MAX5: STD_LOGIC_VECTOR := "100010111101001000"; --143176(DEC)

SIGNAL CONT6 : STD_LOGIC_VECTOR (16 DOWNTO 0) := (OTHERS => '0');
CONSTANT CONT_MAX6: STD_LOGIC_VECTOR := "11000101101110111"; --101239(DEC)

BEGIN
------------------------- PROCESOS DE FRECUENCIAS ---------------------
PROCESS(CLK)
BEGIN
    IF rising_edge(CLK) THEN
        CONT <= CONT + 1;
        IF CONT = CONT_MAX THEN
            CONT <= (OTHERS => '0');
        END IF;

        CONT1 <= CONT1 + 1;
        IF CONT1 = CONT_MAX1 THEN
            CONT1 <= (OTHERS => '0');
        END IF;

        CONT2 <= CONT2 + 1;
        IF CONT2 = CONT_MAX2 THEN
            CONT2 <= (OTHERS => '0');
        END IF;

        CONT3 <= CONT3 + 1;
        IF CONT3 = CONT_MAX3 THEN
            CONT3 <= (OTHERS => '0');
        END IF;

        CONT4 <= CONT4 + 1;
        IF CONT4 = CONT_MAX4 THEN
            CONT4 <= (OTHERS => '0');
        END IF;

        CONT5 <= CONT5 + 1;
        IF CONT5 = CONT_MAX5 THEN
            CONT5 <= (OTHERS => '0');
        END IF;

        CONT6 <= CONT6 + 1;
        IF CONT6 = CONT_MAX6 THEN
            CONT6 <= (OTHERS => '0');
        END IF;
    END IF;
END PROCESS;

------------------------ GENERACIÓN DEL SONIDO ----------------------------
PROCESS(CLK)
BEGIN
    IF rising_edge(CLK) THEN
        IF LA = '0' THEN
            SONIDO <= CONT(16);
        ELSIF DO = '0' THEN
            SONIDO <= CONT1(17);
        ELSIF MI = '0' THEN
            SONIDO <= CONT2(17);
        ELSIF SOL = '0' THEN
            SONIDO <= CONT3(16);
        ELSIF RE = '0' THEN
            SONIDO <= CONT4(17);
        ELSIF FA = '0' THEN
            SONIDO <= CONT5(17);
        ELSIF SI = '0' THEN
            SONIDO <= CONT6(16);
        ELSE
            SONIDO <= '1';
        END IF;
    END IF;
END PROCESS;

END BEHAVIORAL;
