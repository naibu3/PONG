----------------------------------------------------------------------------------
-- Engineer: EFE ACER
-- Project Name: Pong Game
-- Brief: This module is the one that does the painting job. It contains the dynamic
--        position data belonging to different objects, it scans the screen and compares
--        the positions of the cursors with the position data, then it colors the screen
--        in the desired intersections. 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.Constants.all;

entity Sync is
  Port (clock, left, right, start: in std_logic;     
        difficultyControl: in std_logic_vector(1 downto 0);  
        hSync, vSync: out std_logic;
        r, g, b: out std_logic_vector(3 downto 0);
        collision: out std_logic;
        game_started: out std_logic
        );
end Sync;

architecture Behavioral of Sync is
--Defitions of the bitmaps for different images, they will be stored in the ROM 
type BITMAP1 is array (0 to 60) of std_logic_vector(0 to 299);
type BITMAP2 is array (0 to 46) of std_logic_vector(0 to 399);
type BITMAP3 is array (0 to 164) of std_logic_vector(0 to 199);
type BITMAP4 is array (0 to 63) of std_logic_vector(0 to 399);
--Synchronization Signals
signal hPosCurrent, hPosNext: integer range 1 to TOT_H;
signal vPosCurrent, vPosNext: integer range 1 to TOT_V;
--RGB Signals
signal rgbCurrent, rgbNext: std_logic_vector(11 downto 0);
--Intermediate Signals 
signal messageVisible, paddleVisible, ballVisible, frameVisible, paddleAIVisible, result1Visible, result2Visible, logoVisible, gameLabelVisible, borderVisible: boolean;
signal paddleCursor, paddleAICursor: integer range (FP_H + SP_H + BP_H + 1) to (TOT_H - PADDLE_WIDTH):= FP_H + SP_H + BP_H + VIS_H / 2 - (PADDLE_WIDTH + 1) / 2;
signal paddleLeft, paddleRight, paddleAILeft, paddleAIRight: integer range 0 to PRESCALER_PADDLE:= 0;
signal ballCursorX: integer range (FP_H + SP_H + BP_H + 1) to (TOT_H - BALL_SIDE);
signal ballCursorY: integer range (FP_V + SP_V + BP_V + 1) to (TOT_V - BALL_SIDE);
signal ballMovementCounter: integer:= 0;
signal ballMovement: std_logic:= '0';
signal playing: std_logic;
signal newGame, AIWins, playerWins: std_logic;
signal result1, result2: BITMAP1;
signal message: BITMAP2;
signal logo: BITMAP3;
signal gameLabel: BITMAP4;
signal paddleWidth: integer:= PADDLE_WIDTH;

--Component that provides information about the balls position and game logic
component BallController is
    Port (start, move: in std_logic;
          paddleWidth: in integer;
          paddlePos, paddleAIPos: in integer range TOT_H - VIS_H + 1 to TOT_H - PADDLE_WIDTH;
          xPos: out integer range TOT_H - VIS_H + 1 to TOT_H - BALL_SIDE;
          yPos: out integer range TOT_V - VIS_V + 1 to TOT_V;
          newGame, play, AIWon, playerWon: out std_logic;
          ball_collision: out std_logic
          );
end component;
begin
           
    ballControl: BallController 
        port map (start => start,
                  move => ballMovement, 
                  paddleWidth => paddleWidth,
                  paddlePos => paddleCursor, 
                  paddleAIPos => paddleAICursor,
                  xPos => ballCursorX,
                  yPos => ballCursorY,
                  newGame => newGame, 
                  play =>  playing,
                  AIWon => AIWins,
                  playerWon => playerWins,
                  ball_collision => collision);
    --Bitmap assignments for the images  
    -- AI WON          
    result1 <= ("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111",
                "111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111000000010011111111111111111111111",
                "111111111111111111111111111111111111111111111111111110000101111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111100000000000001111111111111111111111",
                "111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111100101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000101111111111111111111111111000000000000000111111111111111111111",
                "111111111111111111111111111111111111111111111111111100000000011111111111111111111111110111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000111111111111111111111111110000000000000011111111111111111111",
                "111111111111111111111111111111111111111111111111111110000000001111111111111111111111010111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000000111111111111111111111111100000000000000001111111111111111111",
                "111111111111111111111111111111111111111111111111111100000000001111111111111111111110010101111111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111111110000000000000001111111111111111111",
                "111111111111111111111111111111111111111111111111111000000000011111111111111111111110000000111111111111111111111111111111010000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000001111111111111111111111110001000000000000000111111111111111111",
                "111111111111111111111111111111111111111111111111111000000001111111111111111111111110000000111111111111111111111111111111010000000111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111000000111111111111111111111111111100000110000000000011111111111111111",
                "111111111111111111110010000000000001111111111111111100000000011111111111111111111110000000111111111111111111111111111111010000000111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111110010000100111111111111111111111111100110000000000000011111111111111111",
                "111111111111111111100000000000000100111111111111111111000000001111111111111111111100000000111111111111111111111111111111010000000111111111111111111111111111111111111111111111111111001010111111111111111111111111111111111111111111111100001000111111111111111111111111101111111100000000011111111111111111",
                "111111111111111111000000000000000000011111111111111111111100011111111111111111111100000000111111111111111111111111111111100000000111111111111111111111001111111111111111111111111111000000011111111111111111111111111111111111111111111111110001111111111111111111111111101111110100000000011111111111111111",
                "111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000111111111111111111111111111111100000000111111111111111111110010000011111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111000110000000011111111111111111",
                "111111111111111110010000000000000000000111111111111111111111111111111111111111111100000000111111111111111111111111111111100000000111111111111111110000000000100000011111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111110110011110100000001111111111111111",
                "111111111111111110000000000000000000000011111111111111111111111111111111111111111100000000111111111111111111111111111111100000000111111111111111110000000000000001001111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111010111110000000001111111111111111",
                "111111111111111110000000000000000000000011111111111111111111111111111111111111111100000000111111111111111111111111111111101000000111111111111111000000000000000000000001111111111110000000011111111111111111111111111111111111111111111111111111111111111111110111011111111100000000000000001111111111111111",
                "111111111111111110000000000000000000000001111111111111110011111111111111111111111101000000111111111111111111111111111111101000000011111111111111000000000000000000000000111111111110000000011111111111111111111111111111111111111111111111111111111111111111111000111111111101110111000000001111111111111111",
                "111111111111111100000000100000000000000000111111111111001011111111111111111111111101000000011111111111111101111111111111101000000011111111111110000000000000000000000000011111111110000000011111111111111111111111111111111111111111111111111111111111110111111100111111111101111110000000001111111111111111",
                "111111111111111100000000000111110100000000111111111110000000111111111111111111111101000000011111111111110101111111111111101000000011111111111110000000000000000000000000001111111110000000001000000000000001111111111111111111111111111111111111111111010111111110011111111101111110000000001111111111111111",
                "111111111111111100000000011111111000000000011111111111000000011111111111111111111101000000011111111111100101011111111111110000000011111111111101000000000000000000000000000111111110000000000000000000000100111111111111111111111111111111111111111110010101001101000111111111111100000000001111111111111111",
                "111111111111111000000000111111111100000000001111111111000000011111111111111111111110000000011111111111100000001111111111110000000011111111111000000000000100000000000000000111111110000000000000000000000000011111111111111111111111111111111111111110000000011101110010111111111000000000001111111111111111",
                "111111111111111000000000111111111101000000001111111111000000011111111111111111111110000000011111111111100000000111111111110000000011111111111000000000000000111000000000000011111110000000010000000000000000001111111111111111111111111111111111111110000000111101111100111111111100000000001111111111111111",
                "111111111111111000000000111111111110000000001111111100000000011111111111111111111110100000011111111111100000000111111111110000000011111111111000000010010011111111000000000011111110000000000000000000000000000111111111111111111111111111111111111110000000110000000100011111111100000000011111111111111111",
                "111111111111111000000001111111111111000000000111111110000000011111111111111111111110100000001111111111000000001111111111110000000011111111110000000000011111111111100000000001111110000000000000000000000000000011111111111111111111111111111111111100000000111011111001111111111000000100011111111111111111",
                "111111111111110000000001111111111111010000000011111110000000011111111111111111111110100000001111111111000000000111111111110000000011111111110000000000111111111111110000000001111110000000000000000000000000000001111111111111111111111111111111111100000000110111111010000110110010000100111111111111111111",
                "111111111111110000000001111111111111010000000011111110000000011111111111111111111110100000001111111111000000000111111111110000000011111111110000000001111111111111110100000000111110000000000000000000000000000000111111111111111111111111111111111101000000100111110111100001111100001000111111111111111111",
                "111111111111110000000011111111111111100000000011111110000000011111111111111111111111000000001111111111000000000111111111110000000011111111110000000011111111111111111000000000111110000000000110000000000000000000111111111111111111111111111111111101000000010111110110010010101111110001111111111111111111",
                "111111111111110000000000000000000000000000000011111110000000011111111111111111111111010000000111111111000000000011111111110000000011111111100000000011111111111111111010000000111110000000001100111111111000000000111111111111111111111111111111111101000000000111101101000100010111111111111111111111111111",
                "111111111111110000000000000000000000000000000011111110000000011111111111111111111111010000000111111111000000000011111111110000000011111111100000000011111111111111111000000000011110000000010001111111111000000000111111111111111111111111111111111101000000000000100100010000000111111111111111111111111111",
                "111111111111110000000000000000000000000000000011111110000000011111111111111111111111010000000111111111000000000011111111110000000011111111100000000111111111111111111100000000011110000000011111111111111100000000011111111111111111111111111111111110000000000000000000100000001111111111111111111111111111",
                "111111111111100000000000000000000000000000000011111110000000011111111111111111111111100000000111111111000000000001111111110000000011111111100000000111111111111111111101000000011110000000011111111111111101000000011111111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
                "111111111111110000000000000000000000000000000011111110000000011111111111111111111111100000000111111111000000000001111111110000000011111111100000000111111111111111111110000000011110000000011111111111111101000000011111111111111111111111111111111111000000000000000000000000111111111111111111111111111111",
                "111111111111110000000000000000000000000000000011111110000000011111111111111111111111101000000111111111000000000000111111110000000011111111100000000111111111111111111110000000011110000000011111111111111100000000011111111111111111111111111111111111100000000000000000000001100111111111111111111111111111",
                "111111111111110000000000000000000000000000000011111110000000011111111111111111111111101000000011111111000000000000001111110000000011111111101000000111111111111111111110000000011110000000011111111111111110000000011111111111111111111111111111111111100000000000000000000011001111111111111111111111111111",
                "111111111111000000000000000000000000000000000011111110000000011111111111111111111111101000000001111111000000000000001111110000000011111111101000000011111111111111111110000000011110000000011111111111111110100000011111111111111111111111111111111111110000000000000000000100011111111111111111111111111111",
                "111111111111110000000000000000000000000000000011111110000000011111111111111111111111101000000001111110000000000000000011110000000011111111101000000011111111111111111110000000011110000000011111111111111100000000011111111111111111111111111111111111110000000000000000011000111111111111111111111111111111",
                "111111111111110000000011111111111111110000000011111110000000011111111111111111111111110000000000111110000000000000000001110000000011111111101000000000111111111111111000000000011110000000011111111111111100000000011111111111111111111111111111111111110000000100000001000011111111111111111111111111111111",
                "111111111111110000000011111111111111110000000011111110000000011111111111111111111111111000000000011110000000000000000001110000000011111111110000000000011111111111111100000000011110000000011111111111111000000000011111111111111111111111111111111111100000000110110000001111111111111111111111111111111111",
                "111111111111110000000011111111111111110000000011111110000000011111111111111111111111111010000000001010000000000000000000110000000011111111110100000000000000000110110001000000011110000000011111111111111000000000011111111111111111111111111111111111100000000111111111111111111111111111111111111111111111",
                "111111111111110100000011111111111111100000000011111110000000011111111111111111111111111100000000000100000000010000000000110000000011111111110000000000000000011000000000000000111110000000011111111111111000000000111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111",
                "111111111111110100000001111111111111100000000011111110000000011111111111111111111111111110000000000000000000011000000000000000000011111111111100000000000000000000000000000000111110000000011111111111110000000000111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111",
                "111111111111110100000001111111111111101000000111111110000000011111111111111111111111111111000000000000000000111100000000000000000011111111111100000000000000000000000000000000111110000000011111111111110000000001111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111",
                "111111111111110100000001111111111111101000000111111110000000011111111111111111111111111111000000000000000000111101000000000000000011111111111111000000000000000000000000001100111110000000011111111111100000000001111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111",
                "111111111111111000000000111111111111101000000111111110100000011111111111111111111111111111110000000000000000111110000000000000000011111111111111110000000000000000000000001001111110000000011111111111100000000001111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111",
                "111111111111111010000000111111111111101000100111111100100000011111111111111111111111111111110100000000000000111110000000000000000011111111111111111000000000000000000000010001111110000000011111111111100000000011111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111",
                "111111111111111010000000111111111111111000100111111110000010011111111111111111111111111111111000000000000001111111100000000000000111111111111111111110000000000000000001100011111110000000011111111111100000000011111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111",
                "111111111111111000000001111111111111111111100111111111100000011111111111111111111111111111111100000000000001111111101000000000100111111111111111111111111000000000001100001111111110100000011111111111000000000111111111111111111111111111111111111110100000001111111111111111111111111111111111111111111111",
                "111111111111111100000001111111111111111111111111111111111110011111111111111111111111111111111111000000000001111111110000000000100111111111111111111111111111111110000001111111111110100000011111111111010000100111111111111111111111111111111111111110100000001111111111111111111111111111111111111111111111",
                "111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111100000010001111111111000000001000111111111111111111111111111111111111111111111111110100000011111111111010001000111111111111111111111111111111111111110000000011111111111111111111111111111111111111111111111",
                "111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111110000000001111111111111111111111111111111111111111111111111110100010011111111111110001001111111111111111111111111111111111111110100010011111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111000111111111111111111111111111111111111111111111111111111100010011111111111111111001111111111111111111111111111111111111101100010011111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111000110011111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"
);          
    -- You WON
    result2 <= ("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111",
                "111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101111111111111111111111111111111111111111",
                "110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001011111111111111111111111111111111111111",
                "111000111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001001111111111111111111111111111111111111",
                "110000011111111111111111111111111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111",
                "110000001111111111111101111111111111111111111111111111111111111111111111111111111100101011111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010000000011111111111111111111111111111111111",
                "111000000111111111111011111111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111110100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111",
                "110000000111111111110100011111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111110100000001111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111",
                "111000000011111111100000001111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111110100000001111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111",
                "111100000011111111100000001111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111110100000001111111111111111111111111111111111111111111111111110010101111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111",
                "111100000001111111000000011111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111000000001111111111111111111110011111111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111",
                "111110000001111111000000011111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111000000001111111111111111111100100000111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111",
                "111110000000111111000000101111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111000000001111111111111111100000000001000000111111111111111110000000111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111",
                "111111000000111110000000011111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111000000001111111111111111100000000000000010011111111111111100000000111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111",
                "111111000000111110000001011111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111010000001111111111111110000000000000000000000011111111111100000000111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111",
                "111111100000011110000000111111111111111111111111111111111111111111111111111111111010000001111111111111111111111111111111010000000111111111111110000000000000000000000001111111111100000000111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111",
                "111111100000001100000000111111111111111111111111111111111111111111111111111111111010000000111111111111111011111111111111010000000111111111111100000000000000000000000000111111111100000000111111111111111111111111111111111111111111111111010111111111110000000000000000000111111111111111111111111111111111",
                "111111100000001100000001111111111111111111111111111111111111111111111111111111111010000000111111111111101011111111111111010000000111111111111100000000000000000000000000011111111100000000010000000000000011111111111111111111111111111100000000000000000000000000000000000011111111111111111111111111111111",
                "111111110000000000000001111111111111111111111111111111111111111111111111111111111010000000111111111111001010111111111111100000000111111111111010000000000000000000000000001111111100000000000000000000001001111111111111111111111111111100000000000000000000000000000000000010101110111111111111111111111111",
                "111111110000000000000001111111111111111111111111110001111111111111111111111111111100000000111111111111000000011111111111100000000111111111110000000000001000000000000000001111111100000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111",
                "111111111000000000000011111111000001111111111111100011111111111111111111111111111100000000111111111111000000001111111111100000000111111111110000000000000001110000000000000111111100000000100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000001111111111111111111",
                "111111111000000000000011111100000010001111111111000000011111111111111111111111111101000000111111111111000000001111111111100000000111111111110000000100100111111110000000000111111100000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000001111111111111111111",
                "111111111100000000001011100001000000001111111111000000001111111111111111111111111101000000011111111110000000011111111111100000000111111111100000000000111111111111000000000011111100000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111",
                "111111111110000000000111100100000000000011111110000000001111111111111111111111111101000000011111111110000000001111111111100000000111111111100000000001111111111111100000000011111100000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111",
                "111111111111000000010110000000000000000001111111000000011111101111111111111111111101000000011111111110000000001111111111100000000111111111100000000011111111111111101000000001111100000000000000000000000000000001111111111111111111101000000000000000000000000000000000000000000000000000000111111111111111",
                "111111111111000000001100100000000000000001111110000001111111000111111111111111111110000000011111111110000000001111111111100000000111111111100000000111111111111111110000000001111100000000001100000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000111111111111111",
                "111111111111000000101000000000000000000000111110000000001110000011111111111111111110100000001111111110000000000111111111100000000111111111000000000111111111111111110100000001111100000000011001111111110000000001111111111111111111111110000000000000000000000000000000000000000000000000000111111111111111",
                "111111111111000000010000000000111000000000011110000000111110000001111111111111111110100000001111111110000000000111111111100000000111111111000000000111111111111111110000000000111100000000100011111111110000000001111111111111111111111111110000000000000000000000000000000000000000000000011111111111111111",
                "111111111110000000000000000001100111000000011111000001111110000000111111111111111110100000001111111110000000000111111111100000000111111111000000001111111111111111111000000000111100000000111111111111111000000000111111111111111111111111111000000000000000000000000000000000000000000001111111111111111111",
                "111111111110000000100000000110011111000000011111000001111110000000111111111111111111000000001111111110000000000011111111100000000111111111000000001111111111111111111010000000111100000000111111111111111010000000111111111111111111111111111100000000000000000000000000000000000000000001111111111111111111",
                "111111111100000000100000001100111111000000011111000000111100000000111111111111111111000000001111111110000000000011111111100000000111111111000000001111111111111111111100000000111100000000111111111111111010000000111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111",
                "111111111100000010100000010011111110000000011111000000000000000000111111111111111111010000001111111110000000000001111111100000000111111111000000001111111111111111111100000000111100000000111111111111111000000000111111111111111111111111111111000000000000000000000000000000000000010000000111111111111111",
                "111111111000000001110000001111111110000000011111000000000010000000111111111111111111010000000111111110000000000000011111100000000111111111010000001111111111111111111100000000111100000000111111111111111100000000111111111111111111111111111110000000000000000000000000000000001110000001111111111111111111",
                "111111111000000101110000000000000000000000011111000000000000000000011111111111111111010000000011111110000000000000011111100000000111111111010000000111111111111111111100000000111100000000111111111111111101000000111111111111111111111111111110000000000000000000000000000000000000000001111111111111111111",
                "111111111000000011110000000000000010000000011111100000000000000000011111111111111111010000000011111100000000000000000111100000000111111111010000000111111111111111111100000000111100000000111111111111111000000000111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111",
                "111111110000001011110000000000000000000000111111100000000000000000011111111111111111100000000001111100000000000000000011100000000111111111010000000001111111111111110000000000111100000000111111111111111000000000111111111111111111111111111100000000000000000000000000000000001111111111111111111111111111",
                "111111110000000111110000000000000000000010111111110000000000010000011111111111111111110000000000111100000000000000000011100000000111111111100000000000111111111111111000000000111100000000111111111111110000000000111111111111111111111111111000000000000000000000000000000000001111111111111111111111111111",
                "111111100000000111111000000000000000001101111111111100000001110000001111111111111111110100000000010100000000000000000001100000000111111111101000000000000000001101100010000000111100000000111111111111110000000000111111111111111111111111111000000000000000000000000000000000001111111111111111111111111111",
                "111111100000001111111000000000000000011001111111111111110000000000001111111111111111111000000000001000000000100000000001100000000111111111100000000000000000110000000000000001111100000000111111111111110000000001111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111",
                "111111100000001111111110000000000001110111111111111111111111110000000111111111111111111100000000000000000000110000000000000000000111111111111000000000000000000000000000000001111100000000111111111111100000000001111111111111111111111111100000000000000000000000000000000000000111111111111111111111111111",
                "111111000000001111111111111000000000001111111111111111111111111000000111111111111111111110000000000000000001111000000000000000000111111111111000000000000000000000000000000001111100000000111111111111100000000011111111111111111111111111000000000000000000000000000000000000000111111111111111111111111111",
                "111111000000011111111111111111111111111111111111111111111111111000000011111111111111111110000000000000000001111010000000000000000111111111111110000000000000000000000000011001111100000000111111111111000000000011111111111111111111111111000000000000000000000000000000000000000111111111111111111111111111",
                "111110000000011111111111111111111111111111111111111111111111111100000011111111111111111111100000000000000001111100000000000000000111111111111111100000000000000000000000010011111100000000111111111111000000000011111111111111111111111110000000000000000000000000000000000000001011111111111111111111111111",
                "111110000001011111111111111111111111111111111111111111111111111100000011111111111111111111101000000000000001111100000000000000000111111111111111110000000000000000000000100011111100000000111111111111000000000111111111111111111111111111000000000000000000001100000000000000000011111111111111111111111111",
                "111110000000111111111111111111111111111111111111111111111111111110000011111111111111111111110000000000000011111111000000000000001111111111111111111100000000000000000011000111111100000000111111111111000000000111111111111111111111111111000000000000000000111100100000000000000111111111111111111111111111",
                "111100000000111111111111111111111111111111111111111111111111111110000001111111111111111111111000000000000011111111010000000001001111111111111111111111110000000000011000011111111101000000111111111110000000001111111111111111111111111110000000000000000001111111000000000000000011111111111111111111111111",
                "111100000001111111111111111111111111111111111111111111111111111110000000111111111111111111111110000000000011111111100000000001001111111111111111111111111111111100000011111111111101000000111111111110100001001111111111111111111111111111100000000000000011111111100000000000000001111111111111111111111111",
                "111000000001111111111111111111111111111111111111111111111111111110000000111111111111111111111111000000100011111111110000000010001111111111111111111111111111111111111111111111111101000000111111111110100010001111111111111111111111111100000000000000000111111111110000000000000001111111111111111111111111",
                "111000000101111111111111111111111111111111111111111111111111111111000001111111111111111111111111110000011111111111111100000000011111111111111111111111111111111111111111111111111101000100111111111111100010011111111111111111111111111110000000000000011111111111111100000000000001111111111111111111111111",
                "111000000011111111111111111111111111111111111111111111111111111111100101111111111111111111111111111111001111111111111111110001111111111111111111111111111111111111111111111111111111000100111111111111111110011111111111111111111111111110110000000001111111111111111110100000000111111111111111111111111111",
                "111000000011111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100110000000011111111111111111111000000000111111111111111111111111111",
                "111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001100011111111111111111111111000000111111111111111111111111111",
                "111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000111111111111111111111111111100001111111111111111111111111",
                "111000010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111110001111111111111111111111111",
                "111001101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"
                );          
	-- NEW GAME
	message <= ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111110011111111111111000000001111111100111111110011111111111111111111111111000000001111111100000000001111111100000000111111110011110011111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111110011111111111111000000001111111100111111110011111111111111111111111111000000001111111100000000001111111100000000111111110011110011111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011000011111111111100000000000011110000111111110000111111111111111111111100000000000011110000000000000011110000000000001111000011000000111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011000011111111111100000000000011110000111111110000111111111111111111111100000000000011110000000000000011110000000000001111000011000000111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111000011000011111111110000001111000000110000111111110000111111111111111111110000001111000000110000001111111111000000111100000011000011000000001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111000011000011111111110000001111000000110000111111110000111111111111111111110000001111000000110000001111111111000000111100000011000011000000001111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111000011000011111111110000111111110000110000001111000000111111111111111111110000111111110000110000111111111111000011111111000011000011000000000011000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111000011000011111111110000111111110000110000001111000000111111111111111111110000111111110000110000111111111111000011111111000011000011000000000011000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011000011111111110000000000000000111100000000000011111111111111111111110000000000000000110000111100000011000000000000000011000011000011000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011000011111111110000000000000000111100000000000011111111111111111111110000000000000000110000111100000011000000000000000011000011000011000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111000011111111110000000000000000111111000000001111111111111111111111110000000000000000110000110000000011000000000000000011000011000011110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111000011111111110000000000000000111111000000001111111111111111111111110000000000000000110000110000000011000000000000000011000011000011110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111000011111111110000111111110000111111111100001111111111111111111111110000111111110000110000111111000011000011111111000011000011000011111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111000011111111110000111111110000111111111100001111111111111111111111110000111111110000110000111111000011000011111111000011000011000011111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111000000111111110000111111110000111111111100001111111111111111111111110000111111110000110000001111000011000011111111000011000011000011111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111000000111111110000111111110000111111111100001111111111111111111111110000111111110000110000001111000011000011111111000011000011000011111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111000000000000110000111111110000111111111100001111111111111111111111110000111111110000110000000000000011000011111111000011000011000011111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111000000000000110000111111110000111111111100001111111111111111111111110000111111110000110000000000000011000011111111000011000011000011111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111110000000011111100111111110011111111111100111111111111111111111111111100111111110011111100000000001111110011111111001111001111110011111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111110000000011111100111111110011111111111100111111111111111111111111111100111111110011111100000000001111110011111111001111001111110011111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111000011100001110000111000011111111111100000000111011110111000011111111111100001110000111011110111000000001110000111000011111111111100000111101111011100000000111000000001110000001110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000010000001000000100000010000001111111111000000000010011110010000001111111111000000100000010001110010000000000100000010000001111111111000000011001111001000000000010000000000100000000100011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110010011001000111100011110001111111111111111100111110011110010001111111111111000111100011110000110011111001111100011110011001111111111001110001001111001111100111111111001111100011000100001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110010011001001111100111110011111111111111111100111110011110010011111111111111001111100111110000010011111001111100111110011001111111111001111001001111001111100111111111001111100111100100000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000010010001000011100000110000011111111111111100111110000000010000111111111111001111100001110010000011111001111100001110010001111111111000000011001111001111100111111111001111100111100100100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000110000011000011110000011000001111111111111100111110000000010000111111111111001111100001110011000011111001111100001110000011111111111001000011001111001111100111111111001111100111100100110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111110000111001111111110011111001111111111111100111110011110010011111111111111001111100111110011100011111001111100111110000111111111111001111001001111001111100111111111001111100111100100111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111110000011000111111100011110001111111111111100111110011110010001111111111111000111100011110011110011111001111100011110000011111111111001110001000110001111100111111111001111100011000100111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111110010001000000100000010000001111111111111100111110011110010000001111111111000000100000010011110011111001111100000010010001111111111000000011000000001111100111111111001111100000000100111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111011001100001110000111000011111111111111101111111011110111000011111111111100001110000111011110111111011111110000111011001111111111100000111100000011111101111111111011111110000001110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"
                );          
    logo <= ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111110101111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000110111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001011111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000101111111111111111111",
                "11111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000111111111111111111",
                "11111111111111111111111111111111111111111100000111111100000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000011111111111111111",
                "11111111111111111111111111111111111111111001111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111000100000000000000000000000000000000000000000000001111111111111111",
                "11111111111111111111111111111111111111100111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111100010000000000000000000000000000000000000000000000000111111111111111",
                "11111111111111111111111111111111111110001111000000111111000000000001000000000001111111111111111111111111111111111111111111111111111001000000000000000000000000000001100000000000000000000111111111111111",
                "11111111111111111111111111111111111101000000000000000000111111111110111111111110001111111111111111111111111111111111111111111111100110000000000000000001100000000000001011000000000000000011111111111111",
                "11111111111111111111111111111111110000000000000000000000001111111111100000001111110111111111111111111111111111111111111111111110001000000000000000011000000001111011110111110000000000000011111111111111",
                "11111111111111111111111111111100000000000000011000000000000111111111001111110000001001111111111111111111111111111111111111111000100000000000110000000011111001111100101111111100000000000010111111111111",
                "11111111111111111111111111110000000000001111111111111000000000111110111111111111110000111111001111111111111111111111111111110010000000000010000011110111110110111111011111111100000000000001111111111111",
                "11111111111111111111111111000000000011111111111111111000000000011110111111111111111111111100000011111111111111111111111111001100000000000100000111111011101111011110101111111011000000000000011111111111",
                "11111111111111111111111110000000001111111111111111111111000000001110011111111111111111111101111011111111111111111111111100010000000000100001110111111101011111100101110011110111100000000000111111111111",
                "11111111111111111111111000000000111111111111111111111111110000000011001111111111111111111110000011111110000111111111111001000000000001000111101011111110111111111001111101101111110000000000001111111111",
                "11111111111111111111100000000011111111111111111111111111111000000001101111111111111111111111111111111111110111111111110010000000000000001111011101111101001111111001111110011111110000000000011111111111",
                "11111111111111111111000000000111111111111111111111111111111100000001100111111111111111111111111111111100110111111111001100000000011000111110111110111011110111110110111111001111111000000000001111111111",
                "11111111111111111110000000011111111111111111111100111111100000000000110011111111111111111111111111111111000111111110010000000001100011001101111111000111111011101111001110110111110100000000001111111111",
                "11111111111111111100000001011111111111111111111101111100010111000000011011111111111111111111111111111111111111111100100000000011001011110011111111100111111101011111110101111011101110000000001111111111",
                "11111111111111111000000110111111111111111111111100110011110111100000001011111111111111111111111111111111111111111001000000001100010011110011111111101011111110111111111011111100011110000000000111111111",
                "11111111111111110000001110111111111111111111111111001111111011110000000011111111111111111111111111111111111111110010000000100001101101101100111111011101111101001111110100111110011110000000000111111111",
                "11111111111111100000011110111111111111111111111111011111111011110000000011111111111111111111111111111111111111100100000001100011011110101111011110111110011011110111101111011110101110000000000111111111",
                "11111111111111000000111101111111111111111111111111011111110011111000000001111111111111111111111111111111111110011000000011001100111111001111100101111111100111111011011111101101110010000000000111111111",
                "11111111111111000001111100111111111111111111111111011111111111111000000000011111111111111111111111111111111100100000001100011100111110110111111011111111100111111100111111110011111100000000000111111111",
                "11111111111110000011111110111111111111111111111111011111111111111100000001100000011111111111111111111111111001000000011000111011011101111011110100111111011011111100111111110001111110000000000111111111",
                "11111111111100000111111110000000111111111111111100111111111111111111000001111111001111111111111111111111110010000000110011010111100011111100101111011110111101111011001111101110111110000000000111111111",
                "11111111111000001111111111111100001111101110000001111111111111111100000001111111101111111111111111111111100100000000100111101111110011111111011111101101111110010111110111011111011100000000000111111111",
                "11111111111000011111111111110011100110001000111111111111111111111100000000000000001111110000111111111111001000000011001111010111101101111110101111110011111111101111111010111111101010000000000111111111",
                "11111111110000011111111111101111110001100011111111111111111111111111000000111111111111100110011111111110010000000110001111011001011110111101110011111001111111010111111101111111110010000000000111111111",
                "11111111110000011111111111101111111111010111111111111111111111111110000001111111111111111001111111111101000000010000110110111110011111001101111101110110011111011011111010111111101100000000001111111111",
                "11111111110000011111111111011111111110111111111111111111111111111110000001111111111111111111111111111000000000110011111001111110011111110011111110101111101110111100110111001111011110000000001111111111",
                "11111111100000011111111111011111111110111111111111111111111111111110000000011111111111111111111111111010000001100101111001111101101111110011111111001111110001111111001111110111011110000000001111111111",
                "11111111000001111111111111111111111100111111111000000001111111111111000001000000111111111111111111110000000011001110110110111011110111101101111110110111111001111111001111111010111110000000001111111111",
                "11111111000001111111111111111111111101111111110000000001111111111110000001111100111111111111111111110000000000011111001111010111111011011110011101111011110110111110110111111101111110000000001011111111",
                "11111111000001111100000011111111111100111111100000000000111111111110000001111001111111111111111111110000000100111111001111101111111100111111101011111100101111001110111011111010111100000000001011111111",
                "11111111000001111000000001111111111101111111100000000000011111111110000001110011111111111111111111100000000001011110110111010111111100111111110111111111011111110101111100110111001010000000001011111111",
                "11111111000001110000000000111111111111111111100000000000001111111111000000000111111111111111111111101000000011101101111010111011111011011111101011111110100111111001111111001111110110000000011011111111",
                "11111110000001100000000000111111111111111111000000000000001111111110000001111111111111111111111111000000000011110011111100111100110111101111011100111101111011110110111111001111101010000000011011111111",
                "11111110000011110000000000011111111111111111000000000000001111111100000001111111111111111111111111000000000111111011111100111111001111110110111111011011111101101111001110110111011100000000011011111111",
                "11111100000011100000000000011111111111111111000000001000001111111100000001111111111111111111111110000000000111110101111011011111101111111001111111100111111110011111110101111000111100000000011011111111",
                "11111100000011100001100000011111111111111111000000100000001111111100000011111111111111111111111110000000000111101110110111101111010111111000111111100111111110101111111011111110111100000000010111111111",
                "11111110000001000000100000011111111111111111110000000000001111111110000011111111111111111111111100000000000111011111001111110110111011110111011111011011111101110111110100111101011000000000011011111111",
                "11111100000001000000000000011111111111111111000000000000011111111100000011111111111111111111111100000000001010111111001111111001111101110111101011011100111011111001101111011011101000000000011011111111",
                "11111111000001000000000000011111111111111111000000000000111111111000000111111111111111111111111100000000011101111110110111111001111110101111110110111111010111111110011111100111110000000000111011111111",
                "11111110000001100000000000011111110000111111100000000000111111111000000111000111111111111111111100000000011010111101111001110110111111011111111001111111101111111110011111101011110000000000110111111111",
                "11111111000000100000000000111111100000011111100000000001111000110000001111011011111111111111111000000000110111001101111110101111011110101111111001111111010111111101100111011100100000000000110111111111",
                "11111110000000110000000000011111000000001111110000000011111000000000001111100011111111111111111000000000001111110011111111011111101101110111110110111110111001111011111010111111000000000001110111111111",
                "11111111100000110000000001111110000000001111111100001111100000000000101111111111111111111111111000000001001111110011111110101111110011111011101111011110111110110111111101111111000000000001110111111111",
                "11111111000000011000000011111100000000000111111111111111111000000001011111111111111111111111110000000001010111101101111110110111110011111101011111101101111111001111111010011110000000000011110111111111",
                "11111111000000011111111111111000001000000011111111111111111000000000001111111111111111111111110000000000111001011110111101111011101101111110111111110011111111101111110111101101000000000011101111111111",
                "11111111100000001111111111111000000000000011111111111111111100000000001111111111111111111111110000000001111110111111011011111101011110111101011111110011111111010011101111110010000000000011101111111111",
                "11111111111000000111111111111000000000000111111111111111111111000000000000000000000000111111110000000011111101011111100111111110111111011011101111101100111110111101011111111000000000000011101111111111",
                "11111111110000000111111111111000001110011111111111111111111111100000000111111111111110011111100000000000111011101111100111111101011111100111110111011111011101111110111111110100000000000111101111111111",
                "11111111111000000011111111111111111111111111111111111111111111110000000001111111111110111111100000000011011011110111011011111011101111100111111010111111101011111101011111101100000000000111011111111111",
                "11111111111100000000000111111111111111111111111111111111111111111000000001000001111110111111100000000111100111111010111101110111110111101011111101111111110111111011100111011000000000001111011111111111",
                "11111111111110000000000111111111111111111111111111110001111111111000000000010010000000111111100000000111100111111101111110101111111011011101111010111111101011111011111010110000000000001111011111111111",
                "11111111111111000000001111111111111111111111111111110001111111111100000011111111111111111111100000000111011011111010011111001111111100111110110111011111011101110111111101110000000000011111011111111111",
                "11111111111111100000001100011111111111111100011111000000111111111000000111111111111111111111100000000000111100110111101111001111111100111111001111101110111110101111111010100000000000011110111111111111",
                "11111111111111100000011000010000111111111100011111000000111111100000000011110001111111111111000000000100111111010111110110110111111011011111001111110101111111011111110111000000000000111110111111111111",
                "11111111111111100000000000110000111111110000011111100000011100000000010000001101111111111111000000000011011111101111111001111011110111101111010111111011111110101111110110000000000000111100111111111111",
                "11111111111111000000000001100001111111110000011111100000011000000001011111110011111111111111000000000111101111010111111001111100101111110110111011110100111101110111101101000000000001111101111111111111",
                "11111111111110000010000011000000111111110000011111110000000000001111000000000111111111111111000000000111110010111011110110111111011111111001111101101111011011111011011000000000000000111101111111111111",
                "11111111111110000000000111000000111111110000001111110000000000111100111111111111111111111111000000000111111101111100101111011110101111111001111110011111100111111100111010000000000000111011111111111111",
                "11111111111100000011000111000001111111110000001111111000000111011001111111111111111111111111000000001001111010111111011111101101110111110110111110011111100111111100010000000000000001111011111111111111",
                "11111111111100000000000111000001111111111000001111111100000011100011111111111111111111111111000000001110110111001110101111110011111011101111011101101111011011111011100000000000000101111011111111111111",
                "11111111111100000000001111000001111111111000000111111110000001101111111111111111111111111111000000001111001111110101110111110101111101011111101011110110111101110111100000000000100101111011111111111111",
                "11111111111000000000011110000011111111111000000111111110000001110111111111111111111111111111000000001111001111111011111001101110111110111111110111111001111110101111000000000001001101110111111111111111",
                "11111111111111000000011110000001111111111100000011111111000000011001111111100111111111111111000000001110110011110101111110101111011101011111110001111001111111001110000000000001001011101111111111111111",
                "11111111111111110000011110000001111111111100000001111111100000011100000000010011111111111110000000001110111101101110011111011111101011101111101110110110111111001100100000000010011011101111111111111111",
                "11111111111111111000011111000001111111111110000000111111110000000111111111110011111111111110000000001101111110011111101110101111110111110111011111001111011110110001000000000000111011101111111111111111",
                "11111111111111111000011111000001111111111110000000011111111000000011111111100111111111111110000000001011111111011111110101110111101011111010111111101111101101110010000000000001110111011111100011111111",
                "11111111111111111000011111000000111111111111100000001111111100000011110000001111111111111100000000000111111110100111111011111001011101111101111111010111110011100100000000000001110111011111001101111111",
                "11111111111111111000011111000000111111111111100000000111111110000011000111111111111111111101000000001111111101111011110100111110011110011010111110111011110011001000000000000011101110111111011101111111",
                "11111111111111111000011111100000111111111111100000000001111110000011011111111111111111111000000000001111111011111101101111011110011111100111011101111101101100010000000000000011101100111110111001111111",
                "11111111111111111000011111100000011111111111110000000000111110000011011111111111111111111000000000000111110111111110011111101101101111100111101011111110011100100000000000000010101101111111000111111111",
                "11111111111111111000001111110000001111111111111100000000001110000011001111111111111111110000000000000111101111111110001111110011110011011011110011111111011001000000000000000001011001111111111111111111",
                "11111111111111111000001111110000000111111111111110000000000100000000011111111111111111110000000000000111011111111101110111110001111100111101101101111110100010000000000000000001011011111111111111111111",
                "11111111111111111000000111111000000111111111111111000000000000001001111111111111111111110000000000000010111111111011111011101110111100111110011110111101100100000000000000000100011011111111111111111111",
                "11111111111111111000000111111100000011111111111111100000000000010011111111111111111111110000000000000011111111110111111100011111011011011110011111011011001000000000000010011100111011111111111111111111",
                "11111111111111111100000011111110000011111111111111100000000000100111111110001111111111100000000000000001111111101111111110011111100111101101100111100110010000001000000100111111110111111111111111111111",
                "11111111111111111100000001111110000000011111111111111000000000011111111101010111111111100000000000000001111111101111111101101111100011110011111011100100100000010000001000110111110111111111111111111111",
                "11111111111111111110000000111111000000011111111111111000000100111111111100110111111111100000000100000000111111011111111011110111011101110101111101010011000000100000001001000011110111111111111111111111",
                "11111111111111111111000000011111000000000111111111111000001001111111111100001111111111000000000000000000011110111111110111111000111110101110111110000000000000000000010010100111110111111111111111111111",
                "11111111111111111111100000001111110000000111111111100000100111100000111111111111111111000000000010000000001101111111101111111100111111001111011110000000000000000001100101100111110111111111111111111111",
                "11111111111111111111100000000111110000000001111111000000011000001100111111111111111111000000000100000000000011111111011111111011011110110111101001000000000000000001001011010111110111111111111111111111",
                "11111111111111111111110000000011110000000000111100000011000111111001111111111111111110000000001110000000000111111111011111111011101110111011110010000000000000000110011011010111101111111111111111111111",
                "11111111111111111111111100000001111100000000000000001111111110000111111111111111111110000000001111000000000011111110111111110111110001111101100100000000000000000100110010010111101111111111111111111111",
                "11111111111111111111111100000000011100000000000000011111100000111111111111111111111110000000001111100000000001111101111111101111111001111110001000000000000000011001100100110111101111111111111111111111",
                "11111111111111111111111110000000000100000000000001111111001111111111111111111111111100000000011111101000000000111011111111011111110110111000000000000000000000100011101011110111101111111111111111111111",
                "11111111111111111111111111100000000000000111100000011000111111111111111111111111111100000000011111110000000000010111111110111111101111000000000000000000000001000111011011110111001111111111111111111111",
                "11111111111111111111111111110000000000010111111111000111111111111111111111111111111100000000011001110000000000000000011101111111011110000000000000000000000110000110010011110111011111111111111111111111",
                "11111111111111111111111111111110000001111111111111111111111111111111111111111111111000000000110101100000000000000001100000000000000000100000000000000000001000110110110111110111011111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000101110101100000000000000000000000000000010000000000000000000000001110100101111110011011111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011110110111000000000000000000000000000000000000000000000001000000110101011111111100111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011100110111100000000000000000000000000000000000000000000000001001110000111111111100111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111100110111110000000000000000000000000000000000000000000000011001110010111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111110101111111000000000000000000000000000000000000000000000110011111101111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111110001111111110000000000000000000000000000000000000010010001011111101111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111100000000000000000000000000000000000000000001000100111011111011111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111110000000000000000000000000000000000000000000000100010011111011111011111111111110001111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111110000000000000000000000000000000000000000000100000000001111111011111011111111111110010111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111110000000000000000100000000000000000000000000000000000000000000010000100001111111111011110111111111111101110111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000010001111111111111011110111111111111100001111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000001000000001110111111111111111011110111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111100010000000000000000000000000000000000000000000000010000000001100011101111111111111111011110111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111000100000000000000000000000000000000000000000011000000011000001111111101111111111111111011110111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111111001000000000000000000000000000000000000000000000011111000111100000000101111111111111111011101111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111100000001000000000000000000000000000000011111001111111111011111111111110110111111111111111011101111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111111000000111100000000000000000000000000010111111110000011110011111111111110110111111111111111011101111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111110001000111100000000000000000000000001111111111111111000110111111111111110110111111111111111011101111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111100010001111100000000000000000000000011111111111111111110111011111111111110111011111111111111011101111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111111000100011111110000000000000000000001111011111111111111110011011111111111110111011111111111110111011111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111110001000011111110000000000000000000011111011111111111111111011011111111111110111011111111111110111011111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111100010000011111110000100000000000001001110111111111111111111011011111111111110110011111111111110011011111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111111000000000011111111000000000000000111101110111111111111111111011011111111111110110111111111111111011011111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111100000001000011111110000000000000001111101110111111111111111111010111111111111110000111111111111111011011111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111111000000011100011111111000000000000011111101101111111111111111111000111111111111111111111111111111111100111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111110000000111100011111111000000000001111111101101111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111100000001111100011111111100000000111111111001101111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111111000000011111100011111111100000001111111111011011111111110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111100000001111111100001111111000000111111111111011011111111110110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111110000000011111111100001111100000001111111111111011011111111100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111100000000111111111100001111000000011111111111111011011111111100110011111111111111111111111111111111111111111001111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111000000001111111111100001110000000111111111111111011011111111101110111111111111111111111111111111111111111111010111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111110000000011111111111100000000000001111111111111111010111111111101101111111111111111111111111111111111111111111100111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111100010000011111000000000000000000111111111111111111000111111111101100111111111111111111111111111111111111111111110111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111100111111111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111110000000000000000000001010000000001111111111111111111111111111111101110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111100000001100011000111111100000000011111111111111111111111111111111101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111000000011100011111111111000000001111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111110000000111100001111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111000000001111100001111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111110000000011111110001111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111100000000111111110001111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111100000000111111110000111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111110000000000111111111000111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111100000001000111111111000110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111000000111000111111111000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111000001111000111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111100000011111000111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111000000111110000011111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111110000000011100000011111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111110000000011100000011111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111100000000011000000011111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111000000000011000000011111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111000000000010000110001110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111000000000000001110000100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111100000000000001111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111000000000000010010000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111000000000000000011100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111100000000000000000100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111100001110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"
); 
    gameLabel <= ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111000001111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111000000000111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111100000000001110001111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111000000000000111111111111111000000001111100000111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000011111111111110000000111111000000001111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000011111111111100000001111111000010000111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000001111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111110000010001111111111111111111111111111100000000000111111111111111111111111111111111111111100000000000001111111111100000111111111000111000111111110000000011111111111111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111",
                "1111111111110000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111111111111111111100000111001111100000011111111111111111110011000000111111111111111111111111111111111111111100000100000000111111111000001111111111000011100011111111000000011111111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111",
                "1111111111000000000011111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000011111111111111111111111111111000001111000000000000001111100000000001110011000000011111111111111111111111111111111111111100000110000000111111110000011111111111100001100000111111100000001111111111111111111111111111111111111111111111111111111111111110000000000011111111111111111111111111",
                "1111111111110000000011111111111111111111111111000000000001111111111111111111110000001111111111111111000000000000000001111111111111111111111111111000000111100000000110001100000000000000010011100000011111111111111111111111111111111111111100000111000000111111110000011111111111110001110000001111110000001111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111",
                "1111111111111000000000111111111111111111100000000000000000000011111111111111100000011111111111111111111111110000000001111110000000000000000000111000000111111111111111001100001111111000000011100000000000000111111111111111111111111111111100000111000000011111100000111111111111110001111100000000110000000111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111",
                "1111111111100000000000011111111111111110000000000000000000000000000011111111000000111111111111100000000011110000000001110000000000000000000000000000000111111111111111001100111111111110000011110000000000000000001111111000000001111111111000001111100000011111100000111111111111110000001111100000011000000111111111111111111100000000000000011111111111111111111111111000000110000000011111111111111111111111",
                "1111111111100000110000011111111111111110000000000000000000000000000000011111000001100000000111000000000001110010000001000000000000000000000000000000000111111111111111001100111111111111111111110000000000000000000111000000000000111111111000001111100000011111100000111111111111111000000001111110001000000111111111111111111000000000000000011111111111111111111111111000001111000000001111111111111111111111",
                "1111111111100000100000000011111111111000000000001111000000000000000000000111000000000000000011001111111000110011000000000000000000000000000000000000000000111111111111001100111111111111111111111000000000000000000100000000000000001111110000011111110000011111000001111111111111111111100000111110001100000011111111111111100000000000000000011111111111111111111111110000011111110000000111111111111111111111",
                "1111111111000001110000000000000000000000000111111111111111100000000000000001000000001111100011001111111000100011000000000000111111111100010000000000000000011111111111001100111111110000111111111100000110000000000000000000000000001111000000011111110000011111000001111111111100011111111000000000001100000011111111111111100000000000000000000111111111111111111111110000011111110000000011111111111111111111",
                "1111111111000001111100000000000000000000001111111111111111111111000000000000000011111111110011001111111100000011000000000111111111111110011111100000000000001111111111001100111111100000001111111000001111111100000000000001100000000000000000100001111000011111000001111111111100000001111110000000011100000011111111111111000000011111110000000111111110000000011111100000111111111000000011111111111111111111",
                "1111111111110000111000000000000000000000111111111111111111111111111000000000000011111111110000001111111100000111000000001111111111111110000111111110000000001111111111000100111111100000001111111000001111111100000000001111110000000000000000000000100000111111000001111111111100000000111111111111111110000011111111111110000001111111111100000111111000000000001111100000111111111100000001111111111111111111",
                "1111111111000000111100110000000000000001111111111111111111111111111110000000000011111111110000001111111100001111000001111111111111111111000001111111100000001111111111000000111111110000001111111000001111111100000001111111111000000000000000000000100000111111000001111111110000000000000111111111111110000011111111111110000011111111111100000011110000000000000111100001111111111110000000111111111111111111",
                "1111111111110000111100111111111111111111111111111111111111111111111111100000000011111111111000111111111111111111000001111111111111111111100000011100010000001111111111100000111111111100111111110000001111111100000111111111111110111000011000110001100000111111000001111111111110000000000011111111111110000011111111111100000111111111111100000011110000000000000011000000000011111000000000111111111111111111",
                "1111111111100000011100011111111111111111111111111111111111111111111111110000000011111111111111111111111111111110000001111111111111111111111100011000000000001111111111111000111111111111111111110000001111111100000111111111111111111111111111110001100000111111000000111111111111100000000001111111100010000011111111111100000111111111111100000001100000010000000011000000000001110000000000011111111111111111",
                "1111111111100000011110000111111111111111111111111111111111111111111111111000000011111111111111111111111111111110000011111111111111111111111110011000000000001111111111111111111111111111111111110000001111111100000111111111111111111111111111100011100000111111000000111111111111111000000001111110000010000000000000000100000000000111111110000001000001111100000011000000110000110011000000001111111111111111",
                "1111111111100000001111000011111111111111111111110001111111111111111111111000000001111111111111000000000000000000000011111111111110001111111110001000111000001111111111111111111111111111111111110000011111111100000111111111111111111111111111000011000001111111111000111111111111111110000001111100001100000000000000000000000000000001111110000001000011111100000000000011111100110011100000001100000000111111",
                "1111111111100000001111110011111111111111111111110001111111111111111111111111000001111111111111000000000000000001001111111111111110000011111111000000111000001111111111111111111111111111111111110000011111111100000111111111111111111111111111000111000001111111100000111111111111111110000001111000111100000000000000000000000111110001100011000000000011111110000000000111111100110011110000000000000000001111",
                "1111111111110000000011110000011111111111111111110000011111111111111111111110000000111111111111000000000000000000001111111111111110000000111111000000111000001111111111111111111111111100000000000000011111111100000111111111111111111111111110001110000001111111100000111111111111111111111111111000111000000000000000000000000111111001100001000000000111111110000000000111111100000011110000000000000000000011",
                "1111111111111000000000111000001111111111111111000000011111111111111111111111000000111111111100000000000000000000000111111111111000000000011111110011111000000000000011111111111110000000000000000000011111111100000111111111111111111111111110001100000001111111100000111111111111111111111111110001111000001111111110000000000011111000100001110000001111111111000000000111111100000111110000000000000000000011",
                "1111111111111000000000000110000111100011111111111000001111111111111111111111000000111111111111111111111110000000000111111111111110000000011111111111111000000000000000111111111110000000000000000000011111111110000000111111111111111111111100010000000011111111100000011111111111111111111111100001110000011111111111100000000011111000100000100000011111111111000000001111111111111111000000000000110000000011",
                "1111111111111100000000000011100100000011111111110000000111110000011111111111100000011111111111111111111111100000000011111111111110000000011111111111111000000000000000111111111000000000000000000000011111111000000000111111111111111111111000000000000011111111100000011111111111111111111111000011100000011111111111110000000001111100100000111000001111111111000000001111111111111110000000000011111100000011",
                "1111111111111100000000000000000000000011111111111110000010000000011111110001100000011111111111111111111111111000000001111111111111100000011111111111111000000000000000111111111000000000000000001111111111111000000000111111111111000000000000000000000111111111111100011111111111111111111110000111000000111111111111111110000000111100010000010000001111111111100000001111111111110000000000011111111110000011",
                "1111111111111110010000000000000000000011111111111110000000000000011111000000111000011111111111111111111111111100000001111111111111111111111111111111111000000000000000111111111000000111111110001111111111111000000000111111111100000000000000000000100111111111110000011111111111111111111000001110000001111111111111111110000000011100000000010000001111111111100000001111111111100000000011111111111110000011",
                "1111111111111110011110000000000000000011111111111100000000000000011111000000110000011111111111111111111111111110000001111111111111111111111111111111111000001111100000111111111000000111111110001111111111100000000111111111111110000000000000000011000111111111110000011111111111111111100000011100000011111111111111111111000000011110000010001000000111111111100000001111111111000000001111111111111110000011",
                "1111111111111110001111100000000000000011111111111110000000000011111110001100010000001111111111111111111111111110000001111111111111111111111111111111111000001111100000111111111000000011111000001111111111111111111111111111111100000000000000001111001111111111110000011111111111111111000001110000000111111111111111111111100000011111111111000000000111111111110000001111111110000000011111111111111110000011",
                "1111111111111111001110000111111000000011111111111111100000111111111110011100010000001111111111111111111111111111000001111111100011111111111111111111111000001111100000111111111100000011111000000111111111111111111111111111111100000110000011111111001111111111111100011111111111111111000110000000001111111111111111111111110000001111111111000000000111111111110000000111111100000011111111111111111110000011",
                "1111111111111111001110000000001000000011111111111111000000111111111110011100011100001111111111111111111111111111000001111111100011111111111111100111111000001111100000111111111100000011111000000111111111111111111111111111111000000111100100000111001111111111110000011111111111111110000000000000011111111111111111111111110000001111111111110000000111111111100000000111111100000111111111111111111100000111",
                "1111111111111111001110000000001000000001111111111111100000011111111110001100011000001111111111111111111111111111000001111111100000111111111000000011111000001111100000111111111110000011111110000111111111111111111111111111111000001111100000000010001111111111110000001111111111111100000000000000111111111111111111111111110000001111111111111000000111111111000111000111111000001111111111111111111100000111",
                "1111111111111111000110011111001000000001111111111111111000011111111110001100011000001111111111110011111111111110000001111110000000000000000000000011111000001111100000111111111110000001111100000111111111111111111111111111110000001111100000100010011111111111111100001111111111111100000000000011111110000000111111111111111000001111111111111100000111111111001100000111110000000000001111111111111100000111",
                "1111111111111111000110011111001001100001111111111111111100011111111110001110001000001111111111110000111111111000000011111111110000000000000000000011111000001111100000111111111110000001111100000111111111111111110011111111111000001111100001110010011111111111110000001111111111110000000000000011111110000000001111111111111110001111111111111111111111111110001100000111110000000000001111111111111100000111",
                "1111111111111111100110011111001001000001111111111111110000011111111110001110001000001111111111110000000000000000000111111111100000000000000000000011111000001111100000111111111111000001111111000111111110000000000001111111110000001111111111100000011111111111111000001111111111110000000111000011111110000000000111111111111000001111111111111111111111111100011111000111110000000000001111111111111000001111",
                "1111111111111111100110011111001001000001111111111111111100001111111000011110001000001111111111110000000000000000001111111111111000000000000001111111110000001111100000111111111110000001111100000111111110000000000001111111111000001111111111100000111111111111111000001111111111110000001110000011111000000000000011111111111000001111111100111111111111111000111100000011111100000000001111111000000000001111",
                "1111111111111111100010011111000001000001111111111111110000001111111000111100011000001111111111100000000000000000000011111111111111100011111111111111100000001111100000111111111111000000111100000111111110000000000001111111111000001111111111100100111111111111111000000111111111111000001100000011111111110000000000111111111000001111111100011111110000011000111100000011111111111111111111100000000000001111",
                "1111111111111111100000011111000011000001111111111111111100001111111001111100011000001111111111110000000000000000000011111111111111100011111111111110000000001111100000111111111111000000111110000111111000000000000001111111111110001111111111100100111111111111111000000111111111111000000100000111111111111100000000111111111000001111111100011111100000000001111111100011111111111111111111000011110000011111",
                "1111111111111111110000111111111111000001111111111111111000001111111001111000110000011111111111111111111111111110000001111111111110000011111111111110001000001111100000111111111111111000011000001111111111100000011111111111111000000111111111100100111111111111111000000111111111111000000100000010001111111110000000111111111100001111111100011111100110000001111110000011111111111111111111000111100000111111",
                "1111111111111111111111111111111111000001111111111111111000001111111000000001100000011111111111111111111111111100000001111111111111100011111111111110011000001111100000111111111111100000011110001111111111100000011111111111111000000111111111000000111111111111111100000111111111110000000100000000000111111111000000111111110000011111110000011111100111111111111110000011111111111111111110001110000000111111",
                "1111111111111111111111111111111111000001111111111111111000001111111000000011100000111111111111111111111111111110000001111111111111100011111111111110011000001111100000111111111111111100011000001111111111100000111111111111111111000111111111001001111111111111111100000111111111110000000000000000000011111111111111111111110000011111110000011111100111111111111110000001111111111111111000001100000001111111",
                "1111111111111111111111111111111111000001111111111111111000001111111111111111000000111111111111111111111111111111000001111111111110000011111111111110011000001111100000111111111111110000011000001111111111100000111111111111111100000111111111001001111111111111111111000111111111100000000010000001110001111111111111111111110000011111110000011111100111111111111100000001111111111111111000111100000011111111",
                "1111111111111111111111110000011111000001111111111111111111111111111111111110000001111111111111111111111111111111000001111111111110000011111111111100010000001111100000111111111111110000011000001111111111100000111111111111111100000111111111001001111111111111111100000111111111000100000010000000111001111111111111111111100000111111110000011111100111111111111110000001111111111111110001111000001111111111",
                "1111111111111111111111110000011111000001111111111111111111111111111111111110000011111111111111111111111111111111000001111111111111000011111111100000010000011111100000111111111111111100011110001111111111100000111111111111111100000111111111000001111111111111111100000111111111000110000011100000011000000000111111111111000000111111110000011111100111111111111110000000111111111111100001100000011111111111",
                "1111111111111111111111100010011111000000111111111111111111111111111111111100000011111111111111111111111111111111000001111111111110000011111110000001110000001111100000111111111111110000001000001111111111000000111111111111111100000111111111000001111111111111111100000111111110001110000011000000001000000000000011111111000000111111110000011111000111111111111100000000111111111111000011000000011111111111",
                "1111111111111111111111100110011111000000111110011100111111111111111111110000000011111111111111111111111111111111000001111111111110000011111110000111110000001111100000111111111111110000001000001111111111100000111111111111111111000111111111000011111111111111111100000111111110011110000011100000000001111110000001111110000000011111110000000110000111111111111000000000001111111111000100000000111111111111",
                "1111111111111111111111100000011111000000001110000000011111111111111111100000000011111111111111111111111111111111000001111111111100000011111100011111110000001111100000111111111111110000001000001111111111100000111111111111111100000111111111100111111111111111111100000111111110011110000011100000000000010001110000000000000000001111110000000000001111111100000000000000000011111111000000000011111111111111",
                "1111111111111111111111110000111111000000000000000000001111111111111110000000000001111111111111111111111111111110000001111111111100000001111100011110000000001111100000111111111111111000001000001111111111100000111111111111111100000111111111111111000001111111111100000011111000011110000011110000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000111111111111111",
                "1111111111111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111100000000000011111111100000000001100100000000000011111100000011111100000000000001000001111111110000001111111111111111100000111111111111110000000111111111111000011100000011100000011111100000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000001111111111111111",
                "1111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000011000000001100000000000111111111111100000000111111111111110001100111111111110000000000000000000000011111111100000000000000000000000010000000000000000000000000000000000000001111110000000000000000001111111111111111111",
                "1111111111111111111111111111111111111000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000011000000000000000000000000001110000000000000111111111111110001100111111111110000000000000000000000111111111110000000000000000000001111000000000000000111100000000000000100011111111000000000000000111111111111111111111",
                "1111111111111111111111111111111111111111111111111000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000001111000000000000000000000000000000000000000001111111111111110000000111111111111000000000000000000000111111111111110000000000001111111111110000000000001111111111111111001100011111111111100000111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011111000000000000000011000000000000011111111111111110000000000000111111111111000000000000000000000000000000000000000011111111111111111000001111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111001000011111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"
                );
    
    game_started <= playing;
    
    --The process involves the next state logic for the variables
    process(clock)
    begin 

        if clock'event and clock = '1' then
        --Producing the clock signal that will occur in the BallController module
            if ballMovementCounter = PRESCALER_BALL then
                ballMovement <= not ballMovement;
                ballMovementCounter <= 0;
            else 
                ballMovementCounter <= ballMovementCounter + 1;
            end if;
            --Button - paddle control
            if playing = '1' then
                if right = '1' and left = '0' then
                    paddleRight <= paddleRight + 1;
                    paddleLeft <= 0;
                elsif left = '1' and right = '0' then
                    paddleLeft <= paddleLeft + 1;
                    paddleRight <= 0;
                else 
                    paddleRight <= 0;
                    paddleLeft <= 0;
                end if;
                --Adjusting the position of the player's paddle according to the specified constant to avoid debouncing
                if paddleRight = (PRESCALER_PADDLE - 5000) and paddleCursor < TOT_H - paddleWidth then
                    paddleCursor <= paddleCursor + 1;
                elsif paddleLeft = (PRESCALER_PADDLE - 5000) and paddleCursor > FP_H + SP_H + BP_H + 1 then
                    paddleCursor <= paddleCursor - 1;
                end if;  
                --The basic A.I algorithm fot the computer to control a paddle, it follows the ball with a little pseudorandom error   
                if ballCursorX >= paddleAICursor + (ballCursorY mod (ballCursorX mod 5)) * ((ballCursorX) mod (ballCursorY mod 5)) + (paddleCursor * paddleAICursor) mod 5 then
                    paddleAIRight <= paddleAIRight + 1;
                    paddleAILeft <= 0;
                elsif ballCursorX <= paddleAICursor - (ballCursorY mod (ballCursorX mod 5)) * ((ballCursorX) mod (ballCursorY mod 5)) - (paddleCursor * paddleAICursor) mod 5 then 
                    paddleAILeft <= paddleAILeft + 1;
                    paddleAIRight <= 0;
                else 
                    paddleAILeft <= 0;
                    paddleAIRight <= 0;
                end if;
                --Adjusting the position of the computer's paddle according to the specified constant to avoid debouncing    
                if paddleAIRight = PRESCALER_PADDLE and paddleAICursor < TOT_H - PADDLE_WIDTH then
                    paddleAICursor <= paddleAICursor + 1;
                elsif paddleAILeft = PRESCALER_PADDLE and paddleAICursor > FP_H + SP_H + BP_H + 1 then
                    paddleAICursor <= paddleAICursor - 1;
                end if;                
            else --The initial positions of the paddles when the game stops
                paddleCursor <= FP_H + SP_H + BP_H + VIS_H / 2 - (PADDLE_WIDTH + 1) / 2;
                paddleAICursor <= FP_H + SP_H + BP_H + VIS_H / 2 - (PADDLE_WIDTH + 1) / 2;
            end if;
            --Register to update the values of the synchronization adn rgb signals
            hPosCurrent <= hPosNext;
            vPosCurrent <= vPosNext;
            rgbCurrent <= rgbNext;
        end if;
    end process;
    
    --Difficulty selection with a multiplexer
    with difficultyControl select paddleWidth <= 
        PADDLE_WIDTH when "00",
        PADDLE_WIDTH_EASY when "01",
        PADDLE_WIDTH_HARD when "10",
        PADDLE_WIDTH when others;  
    --Cursor Position Selections
    result1Visible <= (vPosCurrent >= FP_V + SP_V + BP_V + (VIS_V / 2) - 135) and (vPosCurrent < FP_V + SP_V + BP_V + (VIS_V / 2) - 74) and
                      (hPosCurrent >= FP_H + SP_H + BP_H + (VIS_H / 2) - 150) and (hPosCurrent < FP_H + SP_H + BP_H + (VIS_H / 2) + 150) and
                       result1(vPosCurrent - (FP_V + SP_V + BP_V + (VIS_V / 2) - 135))(hPosCurrent - (FP_H + SP_H + BP_H + (VIS_H / 2) - 150)) 
                       = '0' and AIWins = '1';                  
    result2Visible <= (vPosCurrent >= FP_V + SP_V + BP_V + (VIS_V / 2) - 135) and (vPosCurrent < FP_V + SP_V + BP_V + (VIS_V / 2) - 74) and
                      (hPosCurrent >= FP_H + SP_H + BP_H + (VIS_H / 2) - 150) and (hPosCurrent < FP_H + SP_H + BP_H + (VIS_H / 2) + 150) and
                      result2(vPosCurrent - (FP_V + SP_V + BP_V + (VIS_V / 2) - 135))(hPosCurrent - (FP_H + SP_H + BP_H + (VIS_H / 2) - 150)) 
                      = '0' and playerWins = '1';
    messageVisible <= (vPosCurrent >= FP_V + SP_V + BP_V + (VIS_V / 2) - 50) and (vPosCurrent < FP_V + SP_V + BP_V + (VIS_V / 2) - 3) and
                      (hPosCurrent >= FP_H + SP_H + BP_H + (VIS_H / 2) - 200) and (hPosCurrent < FP_H + SP_H + BP_H + (VIS_H / 2) + 200) and
                       message(vPosCurrent - (FP_V + SP_V + BP_V + (VIS_V / 2) - 50))(hPosCurrent - (FP_H + SP_H + BP_H + (VIS_H / 2) - 200)) 
                       = '0' and newGame = '1';
    logoVisible <= (vPosCurrent >= FP_V + SP_V + BP_V + (VIS_V / 2) + 45) and (vPosCurrent < FP_V + SP_V + BP_V + (VIS_V / 2) + 210) and
                   (hPosCurrent >= FP_H + SP_H + BP_H + (VIS_H / 2) - 100) and (hPosCurrent < FP_H + SP_H + BP_H + (VIS_H / 2) + 100) and
                    logo(vPosCurrent - (FP_V + SP_V + BP_V + (VIS_V / 2) + 45))(hPosCurrent - (FP_H + SP_H + BP_H + (VIS_H / 2) - 100)) 
                    = '0' and newGame = '1';
    gameLabelVisible <= (vPosCurrent >= FP_V + SP_V + BP_V + (VIS_V / 2) - 138) and (vPosCurrent < FP_V + SP_V + BP_V + (VIS_V / 2) - 74) and
                        (hPosCurrent >= FP_H + SP_H + BP_H + (VIS_H / 2) - 200) and (hPosCurrent < FP_H + SP_H + BP_H + (VIS_H / 2) + 200) and
                        gameLabel(vPosCurrent - (FP_V + SP_V + BP_V + (VIS_V / 2) - 138))(hPosCurrent - (FP_H + SP_H + BP_H + (VIS_H / 2) - 200)) 
                        = '0' and AIWins = '0' and playerWins = '0' and newGame = '1';                                                                          
    paddleVisible <= ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 1) and (hPosCurrent > paddleCursor + 8) and (hPosCurrent < paddleCursor + paddleWidth - 8)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 1) and (hPosCurrent > paddleCursor + 7) and (hPosCurrent < paddleCursor + paddleWidth - 7)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 2) and (hPosCurrent > paddleCursor + 6) and (hPosCurrent < paddleCursor + paddleWidth - 6)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 3) and (hPosCurrent > paddleCursor + 5) and (hPosCurrent < paddleCursor + paddleWidth - 5)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 4) and (hPosCurrent > paddleCursor + 4) and (hPosCurrent < paddleCursor + paddleWidth - 4)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 5) and (hPosCurrent > paddleCursor + 3) and (hPosCurrent < paddleCursor + paddleWidth - 3)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 6) and (hPosCurrent > paddleCursor + 2) and (hPosCurrent < paddleCursor + paddleWidth - 2)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 7) and (hPosCurrent > paddleCursor + 1) and (hPosCurrent < paddleCursor + paddleWidth - 1)) or
                     (((vPosCurrent = TOT_V - PADDLE_HEIGHT + 8) or (vPosCurrent = TOT_V - PADDLE_HEIGHT + 9) or (vPosCurrent = TOT_V - PADDLE_HEIGHT + 10)) 
                     and (hPosCurrent > paddleCursor) and (hPosCurrent < paddleCursor + paddleWidth)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 11) and (hPosCurrent > paddleCursor + 1) and (hPosCurrent < paddleCursor + paddleWidth - 1));
    ballVisible <= (((vPosCurrent = ballCursorY) or (vPosCurrent = ballCursorY + BALL_SIDE)) and (hPosCurrent > ballCursorX + 3) and (hPosCurrent <= ballCursorX + 7)) or
                   (((vPosCurrent = ballCursorY + 1) or (vPosCurrent = ballCursorY + BALL_SIDE - 1)) and (hPosCurrent > ballCursorX + 1) and (hPosCurrent <= ballCursorX + 9)) or
                   (((vPosCurrent = ballCursorY + 2) or (vPosCurrent = ballCursorY + BALL_SIDE - 2)
                   or (vPosCurrent = ballCursorY + 3) or (vPosCurrent = ballCursorY + BALL_SIDE - 3)) and (hPosCurrent > ballCursorX) and (hPosCurrent <= ballCursorX + 10)) or
                   ((vPosCurrent > ballCursorY + 2) and (vPosCurrent <= ballCursorY + 7) and (hPosCurrent >= ballCursorX) and (hPosCurrent <= ballCursorX + 11));
    paddleAIVisible <= ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 11) and (hPosCurrent > paddleAICursor + 8) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 8)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 10) and (hPosCurrent > paddleAICursor + 7) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 7)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 9) and (hPosCurrent > paddleAICursor + 6) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 6)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 8) and (hPosCurrent > paddleAICursor + 5) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 5)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 7) and (hPosCurrent > paddleAICursor + 4) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 4)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 6) and (hPosCurrent > paddleAICursor + 3) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 3)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 5) and (hPosCurrent > paddleAICursor + 2) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 2)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 4) and (hPosCurrent > paddleAICursor + 1) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 1)) or
                       (((vPosCurrent = FP_V + SP_V + BP_V + 1 + 3) or (vPosCurrent = FP_V + SP_V + BP_V + 1 + 2) or (vPosCurrent = FP_V + SP_V + BP_V + 1 + 1)) 
                       and (hPosCurrent > paddleAICursor) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1) and (hPosCurrent > paddleAICursor + 1) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 1));                                          
    borderVisible <= (vPosCurrent = FP_V + SP_V + BP_V + (VIS_V / 2) and newGame = '0');
    --Scanning the Pixels
    hPosNext <= hPosCurrent + 1 when hPosCurrent < TOT_H else 1;
    vPosNext <= vPosCurrent + 1 when hPosCurrent = TOT_H and vPosCurrent < TOT_V else
                1 when hPosCurrent = TOT_H and vPosCurrent = TOT_V else vPosCurrent;
	--Color Selection with a multiplexer
    rgbNext <= "001001101110" when paddleVisible else
               "110111011101" when messageVisible else
               "101111110000" when ballVisible else                     
               "110111011101" when frameVisible or borderVisible else
               "100101000100" when paddleAIVisible else
               "100101000100" when result1Visible else
               "000010101110" when result2Visible else
               "001001101110" when gameLabelVisible else
               "001001101110" when logoVisible else
               "000000000000";    
    --Updating the signals that will go to the VGA port
    hSync <= '0' when (hPosCurrent > FP_H) and (hPosCurrent < FP_H + SP_H + 1) else '1';
    vSync <= '0' when (vPosCurrent > FP_V) and (vPosCurrent < FP_V + SP_V + 1) else '1';
    r <= rgbCurrent(11 downto 8);
    g <= rgbCurrent(7 downto 4);
    b <= rgbCurrent(3 downto 0);    
end Behavioral;
